module execution_unit(
  input wire[31:0] oprl,
  input wire[31:0] oprr,
  input wire[31:0] pc,
  input wire[31:0] func_code,

  output wire[31:0] result
);
endmodule